grammar sos:core:files:abstractSyntax;


nonterminal Term with
   pp,
   moduleName,
   tyEnv, constructorEnv,
   type, upSubst, downSubst, finalSubst,
   downVarTypes, upVarTypes,
   headIsConstructor, headConstructorCurrentModule, isVariable,
   errors,
   location;
propagate errors on Term;

--whether the term is headed by a constructor
synthesized attribute headIsConstructor::Boolean;
--whether the term's head is from the current module or is imported
synthesized attribute headConstructorCurrentModule::Boolean;
--whether the term is a variable
synthesized attribute isVariable::Boolean;

abstract production const
top::Term ::= name::QName
{
  top.pp = name.pp;

  name.constructorEnv = top.constructorEnv;

  top.errors <- name.constrErrors;
  top.type = if name.constrFound
             then freshenType(name.constrType)
             else errorType(location=top.location);

  top.upSubst = top.downSubst;

  top.upVarTypes = top.downVarTypes;

  top.headIsConstructor = true;
  top.headConstructorCurrentModule =
      if name.constrFound
      then addQNameBase(top.moduleName, name.base) ==
           name.fullConstrName
      else true; --if not found, just assume it matches
  top.isVariable = false;
}


abstract production var
top::Term ::= name::String
{
  top.pp = name;

  top.upVarTypes =
      if lookup(name, top.downVarTypes).isJust
      then top.downVarTypes
      else (name, top.type)::top.downVarTypes;
  top.type =
      case lookup(name, top.downVarTypes) of
      | just(ty) -> ty
      | nothing() ->
        varType("__var_" ++ name ++ "_" ++ toString(genInt()),
                location=top.location)
      end;

  top.upSubst = top.downSubst;

  top.headIsConstructor = false;
  top.headConstructorCurrentModule = false; --placeholder
  top.isVariable = true;
}


abstract production num
top::Term ::= int::Integer
{
  top.pp = toString(int);

  top.type = intType(location=top.location);

  top.upSubst = top.downSubst;

  top.upVarTypes = top.downVarTypes;

  top.headIsConstructor = false;
  top.headConstructorCurrentModule = false; --placeholder
  top.isVariable = false;
}


abstract production stringConst
top::Term ::= s::String
{
  top.pp = "\"" ++ s ++ "\"";

  top.type = stringType(location=top.location);

  top.upSubst = top.downSubst;

  top.upVarTypes = top.downVarTypes;

  top.headIsConstructor = false;
  top.headConstructorCurrentModule = false; --placeholder
  top.isVariable = false;
}


abstract production appTerm
top::Term ::= constructor::QName args::TermList
{
  top.pp = constructor.pp ++ "(" ++ args.pp_comma ++ ")";

  args.moduleName = top.moduleName;

  constructor.constructorEnv = top.constructorEnv;
  args.tyEnv = top.tyEnv;
  args.constructorEnv = top.constructorEnv;

  top.errors <- constructor.constrErrors;
  top.type = if constructor.constrFound
             then freshenType(constructor.constrType)
             else errorType(location=top.location);

  args.isConclusion = false;
  args.isExtensibleRule = false;
  args.isTranslationRule = false;
  args.expectedPC = nothing();

  args.lastConstructor = constructor;
  args.expectedTypes =
       if constructor.constrFound
       then just(constructor.constrTypeArgs)
       else nothing();
  args.downSubst = top.downSubst;
  top.upSubst = args.upSubst;
  args.finalSubst = top.finalSubst;

  args.downVarTypes = top.downVarTypes;
  top.upVarTypes = args.upVarTypes;

  top.headIsConstructor = true;
  top.headConstructorCurrentModule =
      if constructor.constrFound
      then addQNameBase(top.moduleName, constructor.base) ==
           constructor.fullConstrName
      else true; --if not found, just assume it matches
  top.isVariable = false;
}


abstract production ascriptionTerm
top::Term ::= tm::Term ty::Type
{
  top.pp = "<" ++ tm.pp ++ " : " ++ ty.pp ++ ">";

  tm.moduleName = top.moduleName;

  tm.constructorEnv = top.constructorEnv;
  tm.tyEnv = top.tyEnv;
  ty.tyEnv = top.tyEnv;

  local unify::TypeUnify =
        typeUnify(tm.type, ty, location=top.location);
  tm.downSubst = top.downSubst;
  unify.downSubst = tm.upSubst;
  top.upSubst = unify.upSubst;
  tm.finalSubst = top.finalSubst;

  top.type = ty;

  tm.downVarTypes = top.downVarTypes;
  top.upVarTypes = tm.upVarTypes;

  top.headIsConstructor = tm.headIsConstructor;
  top.headConstructorCurrentModule = tm.headConstructorCurrentModule;
  top.isVariable = tm.isVariable;
}





nonterminal TermList with
   pp_comma, pp_space,
   moduleName,
   tyEnv, constructorEnv,
   types, upSubst, downSubst, finalSubst,
   expectedTypes, lastConstructor,
   downVarTypes, upVarTypes,
   toList<Term>, len,
   expectedPC, isConclusion, isExtensibleRule, isTranslationRule,
   errors,
   location;
propagate errors on TermList;

--When zero, that is the PC
inherited attribute expectedPC::Maybe<Integer>;

abstract production nilTermList
top::TermList ::=
{
  top.pp_comma = "";
  top.pp_space = "";

  top.toList = [];
  top.len = 0;

  top.upSubst = top.downSubst;

  top.errors <-
      case top.expectedTypes of
      | nothing() -> []
      | just(nilTypeList()) -> []
      | just(consTypeList(x, l)) ->
        [errorMessage("Too many arguments to " ++
            top.lastConstructor.pp, location=top.location)]
      end;

  top.types = nilTypeList(location=top.location);

  top.upVarTypes = top.downVarTypes;
}


abstract production consTermList
top::TermList ::= t::Term rest::TermList
{
  top.pp_comma = if rest.pp_comma == ""
                 then t.pp else t.pp ++ ", " ++ rest.pp_comma;
  top.pp_space = if rest.pp_space == ""
                 then t.pp else t.pp ++ " " ++ rest.pp_space;

  t.moduleName = top.moduleName;
  rest.moduleName = top.moduleName;

  t.tyEnv = top.tyEnv;
  t.constructorEnv = top.constructorEnv;
  rest.tyEnv = top.tyEnv;
  rest.constructorEnv = top.constructorEnv;

  top.toList = t::rest.toList;
  top.len = 1 + rest.len;

  t.downSubst = top.downSubst;
  local unifyFirst::TypeUnify =
      case top.expectedTypes of
      | just(consTypeList(ty, l)) ->
        typeUnify(t.type, ty, location=top.location)
             --unify useless as a placeholder
      | _ -> typeUnify(errorType(location=top.location), t.type,
                       location=top.location)
      end;
  rest.downSubst = t.upSubst;
  unifyFirst.downSubst = rest.upSubst;
  top.upSubst = unifyFirst.upSubst;
  t.finalSubst = top.finalSubst;
  rest.finalSubst = top.finalSubst;

  rest.lastConstructor = top.lastConstructor;
  rest.expectedTypes =
       case top.expectedTypes of
       | just(consTypeList(_, l)) -> just(l)
       | _ -> nothing()
       end;
  top.errors <-
      case top.expectedTypes of
      | just(nilTypeList()) ->
        [errorMessage("Too few arguments to " ++
            top.lastConstructor.pp, location=top.location)]
      | _ -> []
      end;

  top.types = consTypeList(t.type, rest.types, location=top.location);

  t.downVarTypes = top.downVarTypes;
  rest.downVarTypes = t.upVarTypes;
  top.upVarTypes = rest.upVarTypes;

  rest.expectedPC = bind(top.expectedPC, \ x::Integer -> just(x - 1));
  rest.isConclusion = top.isConclusion;
  rest.isExtensibleRule = top.isExtensibleRule;
  rest.isTranslationRule = top.isTranslationRule;
  top.errors <-
      if !top.isConclusion
      then []
      else if !top.isExtensibleRule
      then []
      else case top.expectedPC of
           | just(0) ->
             if top.isTranslationRule
             then if t.isVariable then []
                  else [errorMessage("Primary component of " ++
                           "relation " ++ top.lastConstructor.pp ++
                           " in translation rule must be variable;" ++
                           " found " ++ t.pp, location=top.location)]
             else if sameModule(top.moduleName, top.lastConstructor)
                  then [] --initial definition can define anything
                  else if !t.headIsConstructor
                  then [errorMessage("Primary component of " ++
                           "imported relation " ++
                           top.lastConstructor.pp ++
                           " in rule conclusion must be a constructor",
                           location=top.location)]
                  else if !t.headConstructorCurrentModule
                  then [errorMessage("Primary component of " ++
                           "imported relation " ++
                           top.lastConstructor.pp ++
                           " in rule conclusion must be a " ++
                           "constructor introduced in this module",
                           location=top.location)]
                  else [] --PC built by a new constructor
           | _ -> []
           end;
}

