grammar sos:core:main:abstractSyntax;

inherited attribute funEnv::Env<FunctionEnvItem>;

inherited attribute lastFun::QName;
