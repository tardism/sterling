grammar sos:core:concreteDefs:abstractSyntax;

