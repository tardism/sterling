grammar sos:translation:conc:silver;

imports sos:core:common:abstractSyntax;
imports sos:core:concreteDefs:abstractSyntax;

synthesized attribute silverConc<a>::a;
